library verilog;
use verilog.vl_types.all;
entity DFF_32_tb is
end DFF_32_tb;
