library verilog;
use verilog.vl_types.all;
entity key_test_tb is
end key_test_tb;
