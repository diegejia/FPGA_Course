module yindiao
(
 input  [7:0]  hz_sel,
 output reg [19:0] cycle
) ;
  

always @(*)
begin
  case(hz_sel)
     8'h01   : cycle <= 50_000_000/261  ;  
     8'h02   : cycle <= 50_000_000/293  ; 
     8'h03   : cycle <= 50_000_000/329  ;  
     8'h04   : cycle <= 50_000_000/349  ; 
     8'h05   : cycle <= 50_000_000/392  ;  
     8'h06   : cycle <= 50_000_000/440  ;  
     8'h07   : cycle <= 50_000_000/499  ; 
     8'h11   : cycle <= 50_000_000/523  ;  
     8'h12   : cycle <= 50_000_000/587  ;  
     8'h13   : cycle <= 50_000_000/659  ; 
     8'h14   : cycle <= 50_000_000/698  ; 
     8'h15   : cycle <= 50_000_000/784  ;  
     8'h16   : cycle <= 50_000_000/880  ; 
     8'h17   : cycle <= 50_000_000/998  ; 
     8'h21   : cycle <= 50_000_000/1046 ;  
     8'h22   : cycle <= 50_000_000/1174 ; 
     8'h23   : cycle <= 50_000_000/1318 ; 
     8'h24   : cycle <= 50_000_000/1396 ;  
     8'h25   : cycle <= 50_000_000/1568 ;  
     8'h26   : cycle <= 50_000_000/1760 ;  
     8'h27   : cycle <= 50_000_000/1976 ; 
	   8'h31   : cycle <= 50_000_000/2093 ;
	   8'h32   : cycle <= 50_000_000/2349 ; 
	   8'h33   : cycle <= 50_000_000/2637 ; 
	   8'h34   : cycle <= 50_000_000/2794 ; 
	   8'h35   : cycle <= 50_000_000/3136 ; 
	   8'h36   : cycle <= 50_000_000/3520 ;  
 	   8'h37   : cycle <= 50_000_000/3951 ; 
     8'h41   : cycle <= 50_000_000/130 ; 
     8'h42   : cycle <= 50_000_000/146 ;
     8'h43   : cycle <= 50_000_000/165 ;
     8'h44   : cycle <= 50_000_000/175 ;
     8'h45   : cycle <= 50_000_000/196 ;
     8'h46   : cycle <= 50_000_000/220 ;
     8'h47   : cycle <= 50_000_000/250 ; 

     default : cycle <= 20'd0 ;
  endcase
end

endmodule